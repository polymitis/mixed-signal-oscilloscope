library verilog;
use verilog.vl_types.all;
entity PlotSignal is
    generic(
        COLOR_BLACK     : vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        COLOR_RED       : vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        COLOR_GREEN     : vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        COLOR_YELLOW    : vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        COLOR_BLUE      : vl_logic_vector(0 to 11) := (Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        COLOR_FUCHSIA   : vl_logic_vector(0 to 11) := (Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        COLOR_AQUA      : vl_logic_vector(0 to 11) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        COLOR_WHITE     : vl_logic_vector(0 to 11) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        DISP_NCOL       : integer := 160;
        DISP_NROW       : integer := 120;
        GRID_SIDE       : integer := 30;
        GRID_COLOR      : vl_notype;
        DSIG1_COLOR     : vl_notype;
        DSIG2_COLOR     : vl_notype;
        DSIG3_COLOR     : vl_notype;
        DSIG4_COLOR     : vl_notype;
        ASIG1_COLOR     : vl_notype;
        ASIG2_COLOR     : vl_notype;
        TRG_COLOR       : vl_notype;
        MRK_COLOR       : vl_notype;
        TDIV2           : integer := 20;
        TDIV3           : integer := 50;
        TDIV4           : integer := 80;
        TDIV5           : integer := 110;
        TDIV6           : integer := 140;
        ASCL2           : vl_notype;
        ASCL3           : vl_notype;
        ASCL4           : vl_notype;
        DRAW_ASIG_STATE : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        DRAW_DSIG_STATE : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        DRAW_MSIG_STATE : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0)
    );
    port(
        Clock           : in     vl_logic;
        Reset_n         : in     vl_logic;
        X               : out    vl_logic_vector(7 downto 0);
        Y               : out    vl_logic_vector(7 downto 0);
        WR              : out    vl_logic;
        RGB             : out    vl_logic_vector(11 downto 0);
        DISP_VMRK1      : in     vl_logic_vector(8 downto 0);
        DISP_VMRK2      : in     vl_logic_vector(8 downto 0);
        DISP_HMRK1      : in     vl_logic_vector(8 downto 0);
        DISP_HMRK2      : in     vl_logic_vector(8 downto 0);
        INPUT_SELECT    : in     vl_logic_vector(1 downto 0);
        ADC1_RDO_Add    : out    vl_logic_vector(8 downto 0);
        ADC1_RDO_Req    : out    vl_logic;
        ADC1_RDO_Ack    : in     vl_logic;
        ADC1_RDO_Q      : in     vl_logic_vector(13 downto 0);
        ADC1_RDO_Done   : out    vl_logic;
        ADC1_TDiv       : in     vl_logic_vector(0 downto 0);
        ADC1_VDiv       : in     vl_logic_vector(1 downto 0);
        ADC1_VShift     : in     vl_logic_vector(7 downto 0);
        ADC1_TRG_LVL    : in     vl_logic_vector(13 downto 0);
        ADC2_RDO_Add    : out    vl_logic_vector(8 downto 0);
        ADC2_RDO_Req    : out    vl_logic;
        ADC2_RDO_Ack    : in     vl_logic;
        ADC2_RDO_Q      : in     vl_logic_vector(13 downto 0);
        ADC2_RDO_Done   : out    vl_logic;
        ADC2_TDiv       : in     vl_logic_vector(0 downto 0);
        ADC2_VDiv       : in     vl_logic_vector(1 downto 0);
        ADC2_VShift     : in     vl_logic_vector(7 downto 0);
        ADC2_TRG_LVL    : in     vl_logic_vector(13 downto 0);
        DIG1_RDO_Add    : out    vl_logic_vector(8 downto 0);
        DIG1_RDO_Req    : out    vl_logic;
        DIG1_RDO_Ack    : in     vl_logic;
        DIG1_RDO_Q      : in     vl_logic_vector(0 downto 0);
        DIG1_RDO_Done   : out    vl_logic;
        DIG1_TDiv       : in     vl_logic_vector(0 downto 0);
        DIG1_VShift     : in     vl_logic_vector(7 downto 0);
        DIG2_RDO_Add    : out    vl_logic_vector(8 downto 0);
        DIG2_RDO_Req    : out    vl_logic;
        DIG2_RDO_Ack    : in     vl_logic;
        DIG2_RDO_Q      : in     vl_logic_vector(0 downto 0);
        DIG2_RDO_Done   : out    vl_logic;
        DIG2_TDiv       : in     vl_logic_vector(0 downto 0);
        DIG2_VShift     : in     vl_logic_vector(7 downto 0);
        DIG3_RDO_Add    : out    vl_logic_vector(8 downto 0);
        DIG3_RDO_Req    : out    vl_logic;
        DIG3_RDO_Ack    : in     vl_logic;
        DIG3_RDO_Q      : in     vl_logic_vector(0 downto 0);
        DIG3_RDO_Done   : out    vl_logic;
        DIG3_TDiv       : in     vl_logic_vector(0 downto 0);
        DIG3_VShift     : in     vl_logic_vector(7 downto 0);
        DIG4_RDO_Add    : out    vl_logic_vector(8 downto 0);
        DIG4_RDO_Req    : out    vl_logic;
        DIG4_RDO_Ack    : in     vl_logic;
        DIG4_RDO_Q      : in     vl_logic_vector(0 downto 0);
        DIG4_RDO_Done   : out    vl_logic;
        DIG4_TDiv       : in     vl_logic_vector(0 downto 0);
        DIG4_VShift     : in     vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of COLOR_BLACK : constant is 1;
    attribute mti_svvh_generic_type of COLOR_RED : constant is 1;
    attribute mti_svvh_generic_type of COLOR_GREEN : constant is 1;
    attribute mti_svvh_generic_type of COLOR_YELLOW : constant is 1;
    attribute mti_svvh_generic_type of COLOR_BLUE : constant is 1;
    attribute mti_svvh_generic_type of COLOR_FUCHSIA : constant is 1;
    attribute mti_svvh_generic_type of COLOR_AQUA : constant is 1;
    attribute mti_svvh_generic_type of COLOR_WHITE : constant is 1;
    attribute mti_svvh_generic_type of DISP_NCOL : constant is 1;
    attribute mti_svvh_generic_type of DISP_NROW : constant is 1;
    attribute mti_svvh_generic_type of GRID_SIDE : constant is 1;
    attribute mti_svvh_generic_type of GRID_COLOR : constant is 3;
    attribute mti_svvh_generic_type of DSIG1_COLOR : constant is 3;
    attribute mti_svvh_generic_type of DSIG2_COLOR : constant is 3;
    attribute mti_svvh_generic_type of DSIG3_COLOR : constant is 3;
    attribute mti_svvh_generic_type of DSIG4_COLOR : constant is 3;
    attribute mti_svvh_generic_type of ASIG1_COLOR : constant is 3;
    attribute mti_svvh_generic_type of ASIG2_COLOR : constant is 3;
    attribute mti_svvh_generic_type of TRG_COLOR : constant is 3;
    attribute mti_svvh_generic_type of MRK_COLOR : constant is 3;
    attribute mti_svvh_generic_type of TDIV2 : constant is 1;
    attribute mti_svvh_generic_type of TDIV3 : constant is 1;
    attribute mti_svvh_generic_type of TDIV4 : constant is 1;
    attribute mti_svvh_generic_type of TDIV5 : constant is 1;
    attribute mti_svvh_generic_type of TDIV6 : constant is 1;
    attribute mti_svvh_generic_type of ASCL2 : constant is 3;
    attribute mti_svvh_generic_type of ASCL3 : constant is 3;
    attribute mti_svvh_generic_type of ASCL4 : constant is 3;
    attribute mti_svvh_generic_type of DRAW_ASIG_STATE : constant is 1;
    attribute mti_svvh_generic_type of DRAW_DSIG_STATE : constant is 1;
    attribute mti_svvh_generic_type of DRAW_MSIG_STATE : constant is 1;
end PlotSignal;
